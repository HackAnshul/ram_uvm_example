package ram_r_agt_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "ram_defines.svh"
  `include "ram_env_config.svh"

  `include "ram_r_trans.sv"
  `include "ram_r_seqr.sv"

  `include "ram_r_drv.sv"
  `include "ram_r_mon.sv"
  `include "ram_r_agt.sv"

  `include "ram_r_base_seq.sv"

endpackage

